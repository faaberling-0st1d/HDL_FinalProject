/* [Top Module]
 * The top module of all the submodules.
 */

module Top (
);


endmodule