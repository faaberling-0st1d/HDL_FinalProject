module StateEncoder (
    input clk,
    input rst,
    output reg [1:0]
);